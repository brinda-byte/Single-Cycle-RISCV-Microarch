// Design Name: 
// Module Name: andgat
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module andgat(
    input a,
    input b,
    output y
    );
    assign y = a&b;
endmodule
